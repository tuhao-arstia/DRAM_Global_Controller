interface INIT_PHY();

    // Package.sv INPUT FROM PATTERN
    logic rst_n;
    logic clk1;
    logic clk2;
    logic init_ddr_phy_dram_done;

endinterface