////////////////////////////////////////////////////////////////////////
// Project Name: 
// Task Name   : DRAM Frontend Scheduler
// Module Name : frontend_scheduler
// File Name   : frontend_scheduler.sv
// Description : schedule issued commands
////////////////////////////////////////////////////////////////////////

`define B_COUNTER_WIDTH 8
`include "userType_pkg.sv"
`include "define.sv"
`include "FIFO.sv"


module frontend_scheduler(
                          clk,
                          rst_n,
                          something
);

import usertype::*;

input clk;
input rst_n;





// command decoder
logic 


endmodule

